
`include "cpu.v"
`timescale 1ns/1ns
module testbench();
reg clk;
reg reset;
wire [31:0] writedata, dataadr;
wire memwrite;

// instantiate module to be tested
top dut (clk, reset, writedata, dataadr, memwrite);

// initialize test
initial
begin
reset <= 1; # 22; reset <= 0;
end

// clock
always
begin
clk <= 1; # 5; clk <= 0; # 5;
end

initial begin
   $dumpfile("testbench.vcd");
   $dumpvars(0, testbench);
end

// check results
always @ (negedge clk)
begin
   if (memwrite) begin
      if (dataadr == 84 && writedata == 7) begin
          $display ("Simulation succeeded");
             $stop;
                end 
                   else if (dataadr != 80) begin
                       $display ("Simulation failed");
                           $stop;
                       end
                   end
               end
    endmodule
